Library ieee;


--Will complete one day

