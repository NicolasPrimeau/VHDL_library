Library ieee;

